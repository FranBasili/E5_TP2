module LAM(
	input wire clk,
	input wire [31:0] busC,
	
	output wire [31:0] busR,
	output reg writeR		// Indica escritura en registros
);


endmodule